*SI6925DQ  MCE  5-27-97
*20V 3A 0.041ohm Dual Power MOSFET pkg:SMD8B (A:1,4,3)(B:8,5,6)
.SUBCKT SI6925DQ 10 20 40 40
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  18.5M
RS  40  3  2.03M
RG  20  2  44.1
CGS  2  3  560P
EGD 12  0  2  1  1
VFB 14  0  0
FFB  2  1  VFB  1
CGD 13 14  317P
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD  3 10  DSUB
LS  30 40  7.5N
.MODEL DMOS NMOS (LEVEL=3 VMAX=41.7K THETA=80M ETA=2M VTO=0.5 KP=237)
.MODEL DCGD D (CJO=317P VJ=0.6 M=0.68)
.MODEL DSUB D (IS=310N N=1.5 RS=20.6M BV=20 CJO=577P VJ=0.8 M=0.42 TT=50N)
.MODEL DLIM D (IS=100U)
.ENDS 