*SI4980DY  MCE  5-27-97
*80V 4A 0.066ohm Dual Power MOSFET pkg:SMD8A (A:8,2,1)(B:6,4,3)
.SUBCKT SI4980DY 10 20 40 40
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  30.4M
RS  40  3  2.65M
RG  20  2  40.5
CGS  2  3  780P
EGD 12  0  2  1  1
VFB 14  0  0
FFB  2  1  VFB  1
CGD 13 14  290P
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD  3 10  DSUB
LS  30 40  7.5N
.MODEL DMOS NMOS (LEVEL=3 VMAX=167K THETA=80M ETA=2M VTO=2 KP=48.8)
.MODEL DCGD D (CJO=290P VJ=0.6 M=0.68)
.MODEL DSUB D (IS=15.4N N=1.5 RS=67.6M BV=80 CJO=463P VJ=0.8 M=0.42 TT=75N)
.MODEL DLIM D (IS=100U)
.ENDS 