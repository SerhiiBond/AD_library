* 4-Drein 1-Gate 2-Sours
******************************
.SUBCKT 2N7002K 4 1 2
M1   3 1 2 2 NMOS W=26124u L=0.50u
M2   2 1 2 4 PMOS W=26124u L=0.95u
R1   4 3     RTEMP 4.5E-1
CGS  1 2     24E-12
DBD  2 4     DBD
************************************************************
.MODEL  NMOS       NMOS (LEVEL  = 3          TOX    = 7E-8
+ RS     = 4E-1          RD     = 0          NSUB   = 6.2E16
+ KP     = 1E-5          UO     = 650
+ VMAX   = 0             XJ     = 5E-7       KAPPA  = 8E-2
+ ETA    = 1E-4          TPG    = 1
+ IS     = 0             LD     = 0
+ CGSO   = 0             CGDO   = 0          CGBO   = 0
+ NFS    = 0.8E12        DELTA  = 0.1)
************************************************************
.MODEL  PMOS       PMOS (LEVEL  = 3          TOX    = 7E-8
+NSUB    = 2.6E16        TPG    = -1)
************************************************************
.MODEL DBD D (CJO=13E-12 VJ=0.38 M=0.30
+RS=1 FC=0.1 IS=1E-12 TT=4E-8 N=1 BV=60.5)
************************************************************
.MODEL RTEMP RES (TC1=8E-3 TC2=5.5E-6)
************************************************************
.ENDS
