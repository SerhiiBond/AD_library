*BZT52C4V3 MCE 4/8/98
*Ref: Diodes Incorporated, 1994
*4.3V 410mW Si Zener pkg:60A2 1,2
.SUBCKT BZT52C4V3 1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  3.607
.MODEL DF D (IS=2.06N RS=0.102 N=1.7 CJO=100P VJ=0.75 M=0.33 TT=50.1N)
.MODEL DR D (IS=1.02M RS=27 N=12)
.ENDS