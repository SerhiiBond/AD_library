*1N4745A MCE 5/30/96
*Ref: National Discrete Products Databook, 1996
*16V 1W Si pkg:DIODE0.4 1,2
.SUBCKT 1N4745A  1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  15.42
.MODEL DF D (IS=5.02N RS=42M N=1.7 CJO=74.4P VJ=1 M=0.33 TT=50.1N)
.MODEL DR D (IS=870U RS=4.8 N=6.7)
.ENDS 


