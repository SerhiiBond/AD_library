*1N959B MCE 5/30/96
*Ref: National Discrete Products Databook, 1996
*8.2V 500mW Si pkg:DIODE0.4 1,2
.SUBCKT 1N959B   1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  7.671
.MODEL DF D (IS=2.51N RS=84M N=1.7 CJO=46.4P VJ=0.75 M=0.33 TT=50.1N)
.MODEL DR D (IS=9.87U RS=1.95 N=2.6)
.ENDS 


