*DZ23C6V8 MCE 4/9/98
*Ref: Diodes Incorporated, 1994
*6.8V 350mW Si Dual Zener pkg:TO236AA 1,3,2
.SUBCKT DZ23C6V8 1 2 3
*      TERMINALS A K A
XA 1 2 DDZ23C6V8
XB 3 2 DDZ23C6V8
.ENDS DZ23C6V8


.SUBCKT DDZ23C6V8 1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  6.278
.MODEL DF D (IS=1.76N RS=0.12 N=1.7 CJO=43P VJ=0.75 M=0.33 TT=50.1N)
.MODEL DR D (IS=365N RS=4.5 N=2)
.ENDS DDZ23C6V8