*ZPY20 MCE 4/8/98
*Ref: Diodes Incorporated, 1994
*20V 1.3W Si Zener pkg:DIODE0.7 1,2
.SUBCKT ZPY20    1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  19.39
.MODEL DF D (IS=6.53N RS=32.3M N=1.7 CJO=76.8P VJ=1 M=0.33 TT=50.1N)
.MODEL DR D (IS=2.31M RS=3.6 N=8.1)
.ENDS