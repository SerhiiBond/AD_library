*BZT52C12 MCE 4/8/98
*Ref: Diodes Incorporated, 1994
*12V 410mW Si Zener pkg:60A2 1,2
.SUBCKT BZT52C12 1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  11.46
.MODEL DF D (IS=2.06N RS=0.102 N=1.7 CJO=47.5P VJ=1 M=0.33 TT=50.1N)
.MODEL DR D (IS=16.5U RS=7.5 N=3.4)
.ENDS