************ Power Discrete BJT Electrical Parameters ***************
** Product: FJL4215
** Package: TO-264
** Audio Power Amplifier (Complement to FJL4315)
**-------------------------------------------------------------------
.subckt FJL4215 1 2 3
q1 1 2 3 F4215
.model F4215 PNP
+ IS=1.30E-10          BF=91.42             VAF=100
+ IKF=4.480            ISE=1.02E-10         NE=2.0
+ VAR=100              ISC=5.0900E-9        NC=1.5
+ BR=0.882             IKR=2.9015           RE=0.0011
+ RC=0.0553            RB=140.05            RBM=0.0041
+ IRB=8.5e-9           CJE=2.00E-10         FC=0.5
+ CJC=9.45E-10         VJC=0.48             MJC=0.28
+ TF=9.250E-10         XTF=10               VTF=10
+ ITF=1                TR=1.00E-8           EG=0.76
+ XTB=2.68             
.ends FJL4215

***************** Power Discrete Bipolar Thermal Model ****************
.subckt FJL4215_Thermal TH TL
CTHERM1 TH 6 1.84e-3
CTHERM2 6 5  4.24e-3
CTHERM3 5 4  4.62e-3
CTHERM4 4 3  6.24e-3
CTHERM5 3 2  7.02e-2
CTHERM6 2 TL 8.02e-2
RTHERM1 TH 6 2.30e-3
RTHERM2 6 5  1.10e-2
RTHERM3 5 4  1.70e-2
RTHERM4 4 3  2.00e-1
RTHERM5 3 2  2.40e-1
RTHERM6 2 TL 3.50e-1
.ends FJL4315_Thermal 
**-------------------------------------------------------------------
** Creation: Oct.-29-2007   Rev: 1.0
** Fairchild Semiconductor

