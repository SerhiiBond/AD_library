*DZ23C7V5 MCE 4/9/98
*Ref: Diodes Incorporated, 1994
*7.5V 350mW Si Dual Zener pkg:TO236AA 1,3,2
.SUBCKT DZ23C7V5 1 2 3
*      TERMINALS A K A
XA 1 2 DDZ23C7V5
XB 3 2 DDZ23C7V5
.ENDS DZ23C7V5


.SUBCKT DDZ23C7V5 1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  6.978
.MODEL DF D (IS=1.76N RS=0.12 N=1.7 CJO=37.1P VJ=0.75 M=0.33 TT=50.1N)
.MODEL DR D (IS=365N RS=4.5 N=2)
.ENDS DDZ23C7V5