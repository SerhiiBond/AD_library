*1N5358B MCE 6/20/97
*Ref: Diodes Incorporated, 1994
*22V 5W Si Zener pkg:Diode0.7 1,2
.SUBCKT 1N5358B  1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  21.45
.MODEL DF D (IS=5.02N RS=42M N=1.7 CJO=58.2P VJ=1 M=0.33 TT=50.1N)
.MODEL DR D (IS=844U RS=1.05 N=4.7)
.ENDS