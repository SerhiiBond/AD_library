*Si4936DY Siliconix 13-Feb-96
*N-Channel DMOS Subcircuit Model
.SUBCKT Si4936DY 4 1 2 2
M1 3 1 2 2 NMOS W=1232400U L=0.5U
R1 4 3 RTEMP 19M
CGS 1 2 550PF
CGD 1 6 800PF
DMIN 6 4 DMIN
DMAX 6 1 DMAX
DBODY 2 4 DBODY
.MODEL NMOS NMOS(LEVEL=3 TOX=5.0E-8 RS=11M RD=0 LD=0
+ NSUB=1.78E+17 UO=400 VMAX=0 ETA=3.0E-4 XJ=5E-7
+ KAPPA=0 CGBO=0 TPG=1 DELTA=0.1 CGSO=0 CGDO=0
+ IS=0 KP=1.45E-5 NFS=.8E+12)
.MODEL DMIN D(CJO=450E-12 VJ=0.12 M=0.4 FC=0.5 IS=1E-15)
.MODEL DMAX D(CJO=200E-12 VJ=0.8 M=0.5 FC=0.5 IS=1E-15)
.MODEL DBODY D(CJO=840E-12 VJ=0.65 M=0.4 FC=0.5 N=1 IS=1E-15
+ TT=5.7E-8 BV=40)
.MODEL RTEMP R(TC1=7.7M TC2=10U)
.ENDS 