*SUP60N06-18 Siliconix 16-May-96
*N-Channel DMOS Subcircuit Model
.SUBCKT SUP60N06-18 4 1 2 2
M1 3 1 2 2 NMOS W=3525000U L=0.5U
R1 4 3 RTEMP 5M
CGS 1 2 1360PF
CGD 1 6 2000PF
DMIN 6 4 DMIN
DMAX 6 1 DMAX
DBODY 2 4 DBODY
.MODEL NMOS NMOS(LEVEL=3 TOX=80N RS=7M RD=0 LD=0
+ NSUB=4E+15 VTO=4.53 UO=380 VMAX=600K ETA=0.3M XJ=100N THETA=150M
+ KAPPA=0.05 CGBO=0 TPG=1 DELTA=0.1 CGSO=0 CGDO=0 IS=0 NFS=0.5E+10)
.MODEL DMIN D(CJO=1900P VJ=0.08 M=0.58 FC=0.5 IS=1E-20 TT=10N)
.MODEL DMAX D(CJO=900P VJ=0.06 M=0.9 FC=0.5 IS=1E-16 TT=10N)
.MODEL DBODY D(CJO=1350P VJ=0.5 M=0.36 FC=0.5 N=1 IS=1E-15
+ TT=14N BV=68)
.MODEL RTEMP R(TC1=12M TC2=20U)
.ENDS 