*1N4763A MCE 6/20/97
*Ref: Diodes Incorporated, 1994
*91V 1000mW Si Zener pkg:Diode0.7 1,2
.SUBCKT 1N4763A  1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  90.14
.MODEL DF D (IS=5.02N RS=42M N=1.7 CJO=25.4P VJ=1 M=0.33 TT=50.1N)
.MODEL DR D (IS=1.01M RS=75 N=19)
.ENDS