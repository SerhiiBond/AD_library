*DL4730A MCE 4/8/98
*Ref: Diodes Incorporated, 1994
*3.9V 1W Si Zener pkg:DL-41 1,2
.SUBCKT DL4730A  1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  3.125
.MODEL DF D (IS=5.02N RS=42M N=1.7 CJO=283P VJ=0.75 M=0.33 TT=50.1N)
.MODEL DR D (IS=18.5M RS=2.7 N=16)
.ENDS