*DZ23C43 MCE 4/9/98
*Ref: Diodes Incorporated, 1994
*43V 350mW Si Dual Zener pkg:TO236AA 1,3,2
.SUBCKT DZ23C43 1 2 3
*      TERMINALS A K A
XA 1 2 DDZ23C43
XB 3 2 DDZ23C43
.ENDS DZ23C43


.SUBCKT DDZ23C43  1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  42.39
.MODEL DF D (IS=1.76N RS=0.12 N=1.7 CJO=22.7P VJ=1 M=0.33 TT=50.1N)
.MODEL DR D (IS=185U RS=45 N=8.1)
.ENDS DDZ23C43