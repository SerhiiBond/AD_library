*1N5246B MCE 6/2/96
*Ref: National Discrete Products Databook, 1996
*16V 500mW Si pkg:DIODE0.4 1,2
.SUBCKT 1N5246B  1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  15.46
.MODEL DF D (IS=2.51N RS=84M N=1.7 CJO=44.7P VJ=1 M=0.33 TT=50.1N)
.MODEL DR D (IS=35.7U RS=5.1 N=3.6)
.ENDS 


