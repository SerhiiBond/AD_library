*1N5259B MCE 6/20/97
*Ref: Diodes Incorporated, 1994
*39V 500mW Si Zener pkg:Diode0.7 1,2
.SUBCKT 1N5259B  1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  38.41
.MODEL DF D (IS=5.02N RS=42M N=1.7 CJO=39.4P VJ=1 M=0.33 TT=50.1N)
.MODEL DR D (IS=197U RS=24 N=6.9)
.ENDS