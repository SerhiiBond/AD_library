*IRFK3D350 MCE  12/12/97
*Ref: International Rectifier Product Digest '94
*400V 37A .0324ohm Power MOSFET pkg:TO-126 2,3,1
*SYM=POWMOSN
*pn,29/06/2000,merged both parts into 1 subckt

.SUBCKT IRFK3D350 D1 G1 S1D2 G2 S2
X1 D1 G1 S1D2 MIRFK3D350
X2 S1D2 G2 S2 MIRFK3D350
.ENDS

.SUBCKT MIRFK3D350 10 20 40
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  14.4M
RS  40  3  1.81M
RG  20  2  4.05
CGS  2  3  1.07N
EGD 12  0  2  1  1
VFB 14  0  0
FFB  2  1  VFB  1
CGD 13 14  1.35N
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD  3 10  DSUB
LS  30 40  7.5N
.MODEL DMOS NMOS (LEVEL=3 VMAX=833K THETA=58.1M ETA=2M VTO=3.1 KP=10.4)
.MODEL DCGD D (CJO=1.35N VJ=0.6 M=0.68)
.MODEL DSUB D (IS=154N N=1.5 RS=14.9M BV=400 IBV=3M CJO=2.07N VJ=0.8 M=0.42 TT=417N)
.MODEL DLIM D (IS=100U)
.ENDS 
