*ZPY43 MCE 4/8/98
*Ref: Diodes Incorporated, 1994
*43V 1.3W Si Zener pkg:DIODE0.7 1,2
.SUBCKT ZPY43    1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  42.07
.MODEL DF D (IS=6.53N RS=32.3M N=1.7 CJO=43.7P VJ=1 M=0.33 TT=50.1N)
.MODEL DR D (IS=4.09M RS=24 N=22)
.ENDS