*****************************************************************
*SRC=BSS-138;BSS-138;MOSFETs N;Siemens;50V 220mA 3.5 Ohm
*SYM=N-MOSFET
*---------------------------------------------------------------*
* connections:    gate                                          *
*                 | source                                      *
*                 | | drain                                     *
*                 | | |                                         *
.SUBCKT BSS-138   1 2 3
LS 5 2 7N
LD 95 3 5N
RG 4 11 5.5M
RS 5 76 871M
D138 76 95 DREV
.MODEL DREV D CJO=0.06N RS=20M TT=15N IS=300P BV=50
M138 86 11 76 96 MBUZ
.MODEL MBUZ NMOS VTO=1.281 KP=0.186
M2 11 86 8 8 MSW
.MODEL MSW NMOS VTO=0.001 KP=5
M3 86 11 8 8 MSW
COX 11 8 0.08N
DGD 8 86 DCGD
.MODEL DCGD D CJO=0.062N M=0.791 VJ=1.174
CGS 76 11 0.03N
MRDR 86 86 95 86 MVRD
.MODEL MVRD NMOS VTO=-48.9 KP=.045
LG 4 1 7N
.ENDS
