*             G S D
.SUBCKT BSS84 1 2 3
Cgs  2 3 20.6E-12
Cgd1 2 4 56.1E-12
Cgd2 1 4 3.5E-12
M1 1 2 3 3 MOST1 W=12m L=2u
M2 4 2 1 3 MOST2 W=12m L=2u
D1 1 3 Dbody
.MODEL MOST1 PMOS(LEVEL=3 VTO=-1.7 KP=10.07u RD=3.952 RS=20m)
.MODEL MOST2 PMOS(VTO=3.25 KP=10.07u RS=20m)
.MODEL Dbody D(CJO=45.35p VJ=462.4m M=325.5m IS=442f N=1.051 RS=1.243
+              TT=105n BV=50 IBV=10u)
.ENDS
