*BZT52C9V1 MCE 4/8/98
*Ref: Diodes Incorporated, 1994
*9.1V 410mW Si Zener pkg:60A2 1,2
.SUBCKT BZT52C9V1 1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  8.578
.MODEL DF D (IS=2.06N RS=0.102 N=1.7 CJO=32.6P VJ=0.75 M=0.33 TT=50.1N)
.MODEL DR D (IS=365N RS=4.5 N=2)
.ENDS