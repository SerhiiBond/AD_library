*IRFK2F054 MCE  12/12/97
*Ref: International Rectifier Product Digest '94
*60V 120A .01ohm Power MOSFET pkg:TO-126 2,3,1
*SYM=POWMOSN
*pn,27/06/2000,merged both parts into 1 subckt

.SUBCKT IRFK2F054 D1 G1 S1D2 G2 S2
X1 D1 G1 S1D2 MIRFK2F054
X2 S1D2 G2 S2 MIRFK2F054
.ENDS

.SUBCKT MIRFK2F054 10 20 40
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  3.75M
RS  40  3  1.25M
RG  20  2  1.25
CGS  2  3  3.46N
EGD 12  0  2  1  1
VFB 14  0  0
FFB  2  1  VFB  1
CGD 13 14  4.39N
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD  3 10  DSUB
LS  30 40  7.5N
.MODEL DMOS NMOS (LEVEL=3 VMAX=125K THETA=58.1M ETA=2M VTO=3.1 KP=51.6)
.MODEL DCGD D (CJO=4.39N VJ=0.6 M=0.68)
.MODEL DSUB D (IS=498N N=1.5 RS=3.17M BV=60 IBV=2M CJO=6.7N VJ=0.8 M=0.42 TT=593N)
.MODEL DLIM D (IS=100U)
.ENDS 


