*DL5232B MCE 4/8/98
*Ref: Diodes Incorporated, 1994
*5.6V 500mW Si Zener pkg:DL-35 1,2
.SUBCKT DL5232B  1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  5.028
.MODEL DF D (IS=2.51N RS=84M N=1.7 CJO=82.3P VJ=0.75 M=0.33 TT=50.1N)
.MODEL DR D (IS=778U RS=3.3 N=5.9)
.ENDS