*SI3455DV  MCE  5-28-97
* jjt 4/4/2002: changed sign of VTO to match S-56944�Rev. D, 23-Nov-98 datasheet
*30V 4A 0.095ohm Power MOSFET pkg:TSOP-6 1,3,4
.SUBCKT SI3455DV 10 20 40 40
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  44.1M
RS  40  3  3.38M
RG  20  2  42.9
CGS  2  3  410P
EGD 12  0  1  2  1
VFB 14  0  0
FFB  1  2  VFB  1
CGD 13 14  413P
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD 10  3  DSUB
LS  30 40  7.5N
.MODEL DMOS PMOS (LEVEL=3 VMAX=62.5K THETA=80M ETA=2M VTO=-1 KP=8.86)
.MODEL DCGD D (CJO=413P VJ=0.6 M=0.68)
.MODEL DSUB D (IS=14.5N N=1.5 RS=0.129 BV=30 CJO=339P VJ=0.8 M=0.42 TT=50N)
.MODEL DLIM D (IS=100U)
.ENDS 