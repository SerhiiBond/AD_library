*1N5349B MCE 6/20/97
*Ref: Diodes Incorporated, 1994
*12V 5W Si Zener pkg:Diode0.7 1,2
.SUBCKT 1N5349B  1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  11.42
.MODEL DF D (IS=5.02N RS=42M N=1.7 CJO=94.2P VJ=1 M=0.33 TT=50.1N)
.MODEL DR D (IS=5.74M RS=0.75 N=6.8)
.ENDS