*BZT52C22 MCE 4/8/98
*Ref: Diodes Incorporated, 1994
*22V 410mW Si Zener pkg:60A2 1,2
.SUBCKT BZT52C22 1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  21.4
.MODEL DF D (IS=2.06N RS=0.102 N=1.7 CJO=32.7P VJ=1 M=0.33 TT=50.1N)
.MODEL DR D (IS=372U RS=16.5 N=7.4)
.ENDS