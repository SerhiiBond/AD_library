*DZ23C2V7 MCE 4/9/98
*Ref: Diodes Incorporated, 1994
*2.7V 350mW Si Dual Zener pkg:TO236AA 1,3,2
.SUBCKT DZ23C2V7 1 2 3
*      TERMINALS A K A
XA 1 2 DDZ23C2V7
XB 3 2 DDZ23C2V7
.ENDS DZ23C2V7


.SUBCKT DDZ23C2V7 1 2
*     TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  1.975
.MODEL DF D (IS=1.76N RS=0.12 N=1.7 CJO=172P VJ=0.75 M=0.33 TT=50.1N)
.MODEL DR D (IS=1.2M RS=30 N=14)
.ENDS DDZ23C2V7