*IRFK2DE50 MCE  12/12/97
*Ref: International Rectifier Product Digest '94
*800V 12A .1ohm Power MOSFET pkg:TO-126 2,3,1
*SYM=POWMOSN
*pn,27/06/2000,combined subckts into 1 part

.SUBCKT IRFK2DE50 D1 G1 S1D2 G2 S2
X1 D1 G1 S1D2 MIRFK2DE50
X2 S1D2 G2 S2 MIRFK2DE50
.ENDS

.SUBCKT MIRFK2DE50 10 20 40
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  46.5M
RS  40  3  3.5M
RG  20  2  82.5
CGS  2  3  346P
EGD 12  0  2  1  1
VFB 14  0  0
FFB  2  1  VFB  1
CGD 13 14  439P
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD  3 10  DSUB
LS  30 40  7.5N
.MODEL DMOS NMOS (LEVEL=1 LAMBDA=2M VTO=3.1 KP=2.69)
.MODEL DCGD D (CJO=439P VJ=0.6 M=0.68)
.MODEL DSUB D (IS=49.8N N=1.5 RS=62.5M BV=800 IBV=2M CJO=670P VJ=0.8 M=0.42 TT=297N)
.MODEL DLIM D (IS=100U)
.ENDS 


