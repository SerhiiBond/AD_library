*1N4731A MCE 5/30/96
*Ref: National Discrete Products Databook, 1996
*4.3V 1W Si pkg:DIODE0.4 1,2
.SUBCKT 1N4731A  1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  3.561
.MODEL DF D (IS=5.02N RS=42M N=1.7 CJO=244P VJ=0.75 M=0.33 TT=50.1N)
.MODEL DR D (IS=14.8M RS=2.7 N=14)
.ENDS 

