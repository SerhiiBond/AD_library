*DZ23C6V2 MCE 4/9/98
*Ref: Diodes Incorporated, 1994
*6.2V 350mW Si Dual Zener pkg:TO236AA 1,3,2
.SUBCKT DZ23C6V2 1 2 3
*      TERMINALS A K A
XA 1 2 DDZ23C6V2
XB 3 2 DDZ23C6V2
.ENDS DZ23C6V2


.SUBCKT DDZ23C6V2 1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  5.685
.MODEL DF D (IS=1.76N RS=0.12 N=1.7 CJO=49.4P VJ=0.75 M=0.33 TT=50.1N)
.MODEL DR D (IS=3.12N RS=3 N=1.4)
.ENDS DDZ23C6V2