*1N4764A MCE 6/20/97
*Ref: Diodes Incorporated, 1994
*100V 1000mW Si Zener pkg:Diode0.7 1,2
.SUBCKT 1N4764A  1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  99.01
.MODEL DF D (IS=5.02N RS=42M N=1.7 CJO=24.5P VJ=1 M=0.33 TT=50.1N)
.MODEL DR D (IS=1.11M RS=105 N=24)
.ENDS