*DL4753A MCE 4/8/98
*Ref: Diodes Incorporated, 1994
*36V 1W Si Zener pkg:DL-41 1,2
.SUBCKT DL4753A  1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  35.37
.MODEL DF D (IS=5.02N RS=42M N=1.7 CJO=41.4P VJ=1 M=0.33 TT=50.1N)
.MODEL DR D (IS=909U RS=15 N=9.5)
.ENDS