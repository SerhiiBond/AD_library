*ZY130 MCE 4/9/98
*Ref: Diodes Incorporated, 1994
*130V 2W Si Zener pkg:DIODE0.7 1,2
.SUBCKT ZY130    1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  128.5
.MODEL DF D (IS=10N RS=21M N=1.7 CJO=29.6P VJ=1 M=0.33 TT=50.1N)
.MODEL DR D (IS=3.11M RS=90 N=41)
.ENDS