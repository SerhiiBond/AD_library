*Si3441DV Siliconix 21-Oct-96
*P-Channel DMOS Subcircuit Model
.SUBCKT Si3441DV 4 1 2 2
M1 3 1 2 2 PMOS W=300454U L=0.5U
R1 4 3 RTEMP 52.8530M
CGS 1 2 250PF
CGD 1 6 245PF
DMIN 4 6 DMIN
DMAX 1 6 DMAX
DBODY 4 2 DBODY
.MODEL PMOS PMOS(LEVEL=3 TOX=1.75E-8 RS=0.001 RD=0 LD=0
+ NSUB=3.3617E+17 VTO=-1.1738 UO=250 VMAX=0 ETA=3E-4 XJ=0.5E-6
+ KAPPA=0.012 CGBO=0 THETA=0.0 TPG=-1 DELTA=0.0 CGSO=0 CGDO=0
+ IS=0 KP=18.4008U)
.MODEL DMIN D(CJO=1850E-12 VJ=0.12 M=0.72 FC=0.56 IS=1E-20)
.MODEL DMAX D(CJO=1700E-12 VJ=0.50 M=0.5 FC=0.5 IS=1E-22)
.MODEL DBODY D(CJO=420E-12 VJ=0.11 M=0.23 FC=0.5 N=1 IS=1E-18
+ TT=1.0E-7 BV=40)
.MODEL RTEMP R(TC1=4.0E-3 TC2=6.0E-6)
.ENDS Si3441DV