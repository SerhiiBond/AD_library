*DL4761A MCE 4/8/98
*Ref: Diodes Incorporated, 1994
*75V 1W Si Zener pkg:DL-41 1,2
.SUBCKT DL4761A  1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  74.22
.MODEL DF D (IS=5.02N RS=42M N=1.7 CJO=27.7P VJ=1 M=0.33 TT=50.1N)
.MODEL DR D (IS=958U RS=52.5 N=16)
.ENDS