*DL5255B MCE 4/8/98
*Ref: Diodes Incorporated, 1994
*28V 500mW Si Zener pkg:DL-35 1,2
.SUBCKT DL5255B  1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  27.44
.MODEL DF D (IS=2.51N RS=84M N=1.7 CJO=32P VJ=1 M=0.33 TT=50.1N)
.MODEL DR D (IS=122U RS=13.2 N=5.3)
.ENDS