*ZY110 MCE 4/9/98
*Ref: Diodes Incorporated, 1994
*110V 2W Si Zener pkg:DIODE0.7 1,2
.SUBCKT ZY110    1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  108.7
.MODEL DF D (IS=10N RS=21M N=1.7 CJO=32.3P VJ=1 M=0.33 TT=50.1N)
.MODEL DR D (IS=2.82M RS=75 N=34)
.ENDS