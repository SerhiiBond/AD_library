*1N5238B MCE 6/2/96
*Ref: National Discrete Products Databook, 1996
*8.7V 500mW Si pkg:DIODE0.4 1,2
.SUBCKT 1N5238B  1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  8.151
.MODEL DF D (IS=2.51N RS=84M N=1.7 CJO=42.5P VJ=0.75 M=0.33 TT=50.1N)
.MODEL DR D (IS=230U RS=2.4 N=4.3)
.ENDS 


