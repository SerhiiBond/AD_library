*1N749A MCE 5/30/96
*Ref: National Discrete Products Databook, 1996
*4.3V 500mW Si pkg:DIODE0.4 1,2
.SUBCKT 1N749A   1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  3.613
.MODEL DF D (IS=2.51N RS=84M N=1.7 CJO=122P VJ=0.75 M=0.33 TT=50.1N)
.MODEL DR D (IS=3.94M RS=6.6 N=12)
.ENDS 


