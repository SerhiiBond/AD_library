*1N4758A MCE 6/20/97
*Ref: Diodes Incorporated, 1994
*56V 1000mW Si Zener pkg:Diode0.7 1,2
.SUBCKT 1N4758A  1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  55.28
.MODEL DF D (IS=5.02N RS=42M N=1.7 CJO=32P VJ=1 M=0.33 TT=50.1N)
.MODEL DR D (IS=1.06M RS=33 N=13)
.ENDS