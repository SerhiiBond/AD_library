*1N5260B MCE 6/20/97
*Ref: Diodes Incorporated, 1994
*43V 500mW Si Zener pkg:Diode0.7 1,2
.SUBCKT 1N5260B  1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  42.4
.MODEL DF D (IS=5.02N RS=42M N=1.7 CJO=37.1P VJ=1 M=0.33 TT=50.1N)
.MODEL DR D (IS=232U RS=27.9 N=7.5)
.ENDS