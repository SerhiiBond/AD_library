*****************************************************************
*SRC=BSS-92;BSS-92;MOSFETs P;Siemens;240V 150mA 20 Ohm
*SYM=P-MOSFET
 connections:    gate                                           *
*                 | source                                      *
*                 | | drain                                     *
*                 | | |                                         *
.SUBCKT BSS-92    1 2 3
LS 5 2 7N
LD 97 3 5N
RG 86 87 5.5M
RS 5 76 886M
D92 97 76 DREV
.MODEL DREV D CJO=0.05N RS=20M TT=35N IS=300P BV=240
M92 98 87 76 76 MBUZ
.MODEL MBUZ PMOS VTO=-1.489 KP=0.049
M2 87 98 8 8 MSW
.MODEL MSW PMOS VTO=-0.001 KP=5
M3 98 87 8 8 MSW
COX 87 8 0.15N
DGD 98 8 DCGD
.MODEL DCGD D CJO=120P M=0601 VJ=0.47
CGS 76 87 0.06N
MHELP 98 98 97 98 MVRD
.MODEL MVRD PMOS VTO=20.07 KP=0.008
LG 86 1 7N
.ENDS
