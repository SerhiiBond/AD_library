*1N973B MCE 5/30/96
*Ref: National Discrete Products Databook, 1996
*33V 500mW Si pkg:DIODE0.4 1,2
.SUBCKT 1N973B   1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  32.43
.MODEL DF D (IS=2.51N RS=84M N=1.7 CJO=29.4P VJ=1 M=0.33 TT=50.1N)
.MODEL DR D (IS=149U RS=17.4 N=6)
.ENDS 

