*1N754A MCE 5/30/96
*Ref: National Discrete Products Databook, 1996
*6.8V 500mW Si pkg:DIODE0.4 1,2
.SUBCKT 1N754A   1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  6.27
.MODEL DF D (IS=2.51N RS=84M N=1.7 CJO=61.5P VJ=0.75 M=0.33 TT=50.1N)
.MODEL DR D (IS=15.8U RS=1.5 N=2.7)
.ENDS 


