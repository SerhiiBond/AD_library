*ZMU150 MCE 4/8/98
*Ref: Diodes Incorporated, 1994
*150V 1W Si Zener pkg:DL-41 1,2
.SUBCKT ZMU150   1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  148.3
.MODEL DF D (IS=5.02N RS=42M N=1.7 CJO=21.3P VJ=1 M=0.33 TT=50.1N)
.MODEL DR D (IS=3.36M RS=108 N=49)
.ENDS