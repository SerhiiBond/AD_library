*IRGBF30F  MCE  C G E  7-13-95
*900V 20A 17.2ns pkg:TO-220 2,1,3
.SUBCKT IRGBF30F 71 72 74
Q1  83 81 85     QOUT
M1  81 82 83 83  MFIN L=1U W=1U
DSD 83 81  DO
DBE 85 81  DE
RC  85 71  57.2M
RE  83 73  5.72M
RG  72 82  40.2
CGE 82 83  711P
CGC 82 71  1P
EGD 91  0 82 81  1
VFB 93  0  0
FFB 82 81  VFB  1
CGD 92 93  705P
R1  92  0  1
D1  91 92  DLIM
DHV 94 93  DR
R2  91 94  1
D2  94  0  DLIM
LE  73 74  7.5N
DLV 94 95  DR 13
RLV 95  0  1
ESD 96 93  POLY(1) 83 81  19  1
MLV 95 96 93 93  SW
.MODEL SW NMOS (LEVEL=3 VTO=0 KP=5)
.MODEL QOUT PNP (IS=6.23F NF=1.2 BF=5.1 CJE=1.73N TF=17.2N XTB=1.3)
.MODEL MFIN NMOS (LEVEL=3 VMAX=552K THETA=46.1M ETA=1.33M VTO=5.2 KP=1)
.MODEL DR D (IS=.623F CJO=50.3P VJ=1 M=.82)
.MODEL DO D (IS=.623F BV=900 CJO=1.03N VJ=1 M=.7)
.MODEL DE D (IS=.623F BV=14.3 N=2)
.MODEL DLIM D (IS=100N)
.ENDS IRGBF30F 

* Origin: Mceigbts.lib
