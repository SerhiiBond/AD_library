*Si9936DY Siliconix 15-Feb-96
*N-Channel DMOS Subcircuit Model
.SUBCKT Si9936DY 4 1 2 2
M1 3 1 2 2 NMOS W=2453000U L=0.5U
R1 4 3 RTEMP 9.2M
CGS 1 2 80PF
CGD 1 6 900PF
DMIN 6 4 DMIN
DMAX 6 1 DMAX
DBODY 2 4 DBODY
.MODEL NMOS NMOS(LEVEL=3 TOX=50N RS=26M RD=0 LD=0 KP=1.65U
+ NSUB=31.5E+16 UO=500 VMAX=40MEG ETA=0.1M XJ=500N THETA=5M
+ KAPPA=0.08 CGBO=0 TPG=1 DELTA=0.1 CGSO=0 CGDO=0 IS=0 NFS=3E+12)
.MODEL DMIN D(CJO=700P VJ=0.2 M=0.6 FC=0.5)
.MODEL DMAX D(CJO=800P VJ=0.98 M=0.5 FC=0.5 IS=0.5E-15)
.MODEL DBODY D(CJO=900P VJ=0.4 M=0.3 FC=0.5 N=1 IS=1E-10
+ TT=45N BV=40)
.MODEL RTEMP R(TC1=13.5M TC2=50U)
.ENDS 