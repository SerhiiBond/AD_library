*IRGAC50U  MCE  C G E  4/2/98
*Ref: IR Power Semiconductors Product Digest '94
*600V 41A 24.7ns pkg:TO-3 3,2,1
.SUBCKT IRGAC50U 71 72 74
*     TERMINALS:  C  G  E
Q1  83 81 85     QOUT OFF
M1  81 82 83 83  MFIN L=1U W=1U
DSD 83 81  DO
DBE 85 81  DE
RC  85 71  30.2M
RE  83 73  3.02M
RG  72 82  9.76
CGE 82 83  1.88N
EGD 91  0 82 81  1
VFB 93  0  0
FFB 82 81  VFB  1
CGD 92 93  2.09N
R1  92  0  1
D1  91 92  DLIM
DHV 94 93  DR
R2  91 94  1
D2  94  0  DLIM
LE  73 74  7.5N
DLV 94 95  DR 13
RLV 95  0  1
ESD 96 93  POLY(1) 83 81 19  1
MLV 95 96 93 93  SW
.MODEL SW NMOS (LEVEL=3 VTO=0 KP=5)
.MODEL QOUT PNP (IS=387F NF=1.2 BF=5.1 CJE=4.83N TF=24.7N XTB=1.3)
.MODEL MFIN NMOS (LEVEL=3 VMAX=400K THETA=60M ETA=2.01M VTO=4 KP=2.24)
.MODEL DR D (IS=38.7F CJO=149P VJ=1 M=0.82)
.MODEL DO D (IS=38.7F BV=599 CJO=2.74N VJ=1 M=0.7)
.MODEL DE D (IS=38.7F BV=15 N=2)
.MODEL DLIM D (IS=100N)
.ENDS


