*1N5362B MCE 6/20/97
*Ref: Diodes Incorporated, 1994
*28V 5W Si Zener pkg:Diode0.7 1,2
.SUBCKT 1N5362B  1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  27.39
.MODEL DF D (IS=5.02N RS=42M N=1.7 CJO=48.9P VJ=1 M=0.33 TT=50.1N)
.MODEL DR D (IS=4.62M RS=1.8 N=8.1)
.ENDS