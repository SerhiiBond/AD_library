*Si6943DQ Siliconix 01-Aug-95
* jjt 4/4/2002: changed VTO to -0.6V to match S-49534�Rev. E, 06-Oct-97 datasheet.
*P-Channel DMOS Subcircuit Model
.SUBCKT Si6943DQ 4 1 2 2
M1 3 1 2 2 PMOS W=298454U L=0.5U
R1 4 3 RTEMP 8M
CGS 1 2 98PF
CGD 1 6 1195PF
DMIN 4 6 DMIN
DMAX 1 6 DMAX
DBODY 4 2 DBODY
.MODEL PMOS PMOS(LEVEL=3 TOX=17.5N RS=22M RD=0 LD=0 NFS=0.8E+12
+ NSUB=1E+16 UO=400 VTO=-0.6 VMAX=0 ETA=100U XJ=500N
+ KAPPA=1M CGBO=0 TPG=-1 DELTA=0.1 CGSO=0 CGDO=0
+ IS=0 KP=25U)
.MODEL DMIN D(CJO=1617P VJ=0.1 M=0.58 FC=0.5 IS=1E-18)
.MODEL DMAX D(CJO=900P VJ=0.8 M=0.4 FC=0.5 IS=1E-20)
.MODEL DBODY D(CJO=580P VJ=0.15 M=0.26 FC=0.5 N=1 IS=1E-15
+ TT=14N BV=40)
.MODEL RTEMP R(TC1=3.2M TC2=12U)
.ENDS Si6943DQ