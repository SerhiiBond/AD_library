*ZPY4_7 MCE 4/8/98
*Ref: Diodes Incorporated, 1994
*4.7V 1.3W Si Zener pkg:DIODE0.7 1,2
.SUBCKT ZPY4_7   1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  3.839
.MODEL DF D (IS=6.53N RS=32.3M N=1.7 CJO=278P VJ=0.75 M=0.33 TT=50.1N)
.MODEL DR D (IS=36M RS=2.1 N=19)
.ENDS