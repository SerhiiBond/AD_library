*1N5256B MCE 6/2/96
*Ref: National Discrete Products Databook, 1996
*30V 500mW Si pkg:DIODE0.4 1,2
.SUBCKT 1N5256B  1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  29.43
.MODEL DF D (IS=2.51N RS=84M N=1.7 CJO=30.8P VJ=1 M=0.33 TT=50.1N)
.MODEL DR D (IS=131U RS=14.7 N=5.6)
.ENDS 


