*DL5242B MCE 4/8/98
*Ref: Diodes Incorporated, 1994
*12V 500mW Si Zener pkg:DL-35 1,2
.SUBCKT DL5242B  1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  11.21
.MODEL DF D (IS=2.51N RS=84M N=1.7 CJO=54.6P VJ=1 M=0.33 TT=50.1N)
.MODEL DR D (IS=6.08M RS=9 N=16)
.ENDS