*DZ23C24 MCE 4/9/98
*Ref: Diodes Incorporated, 1994
*24V 350mW Si Dual Zener pkg:TO236AA 1,3,2
.SUBCKT DZ23C24 1 2 3
*      TERMINALS A K A
XA 1 2 DDZ23C24
XB 3 2 DDZ23C24
.ENDS DZ23C24


.SUBCKT DDZ23C24  1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  23.37
.MODEL DF D (IS=1.76N RS=0.12 N=1.7 CJO=28.9P VJ=1 M=0.33 TT=50.1N)
.MODEL DR D (IS=650U RS=21 N=9.5)
.ENDS DDZ23C24