*IRGPC50K  MCE  C G E  7-13-95
*600V 55A 28.5ns pkg:TO-247 2,1,3
.SUBCKT IRGPC50K 71 72 74
Q1  83 81 85     QOUT
M1  81 82 83 83  MFIN L=1U W=1U
DSD 83 81  DO
DBE 85 81  DE
RC  85 71  11.5M
RE  83 73  1.15M
RG  72 82  20.3
CGE 82 83  1.95N
CGC 82 71  1P
EGD 91  0 82 81  1
VFB 93  0  0
FFB 82 81  VFB  1
CGD 92 93  1.93N
R1  92  0  1
D1  91 92  DLIM
DHV 94 93  DR
R2  91 94  1
D2  94  0  DLIM
LE  73 74  7.5N
DLV 94 95  DR 13
RLV 95  0  1
ESD 96 93  POLY(1) 83 81  19  1
MLV 95 96 93 93  SW
.MODEL SW NMOS (LEVEL=3 VTO=0 KP=5)
.MODEL QOUT PNP (IS=5.94P NF=1.2 BF=5.1 CJE=4.79N TF=28.5N XTB=1.3)
.MODEL MFIN NMOS (LEVEL=3 VMAX=400K THETA=46.1M ETA=2M VTO=5.2 KP=2.91)
.MODEL DR D (IS=594F CJO=138P VJ=1 M=.82)
.MODEL DO D (IS=594F BV=600 CJO=2.85N VJ=1 M=.7)
.MODEL DE D (IS=594F BV=14.3 N=2)
.MODEL DLIM D (IS=100N)
.ENDS IRGPC50K 


