*******************************************************************
.SUBCKT BDX33B 1 2 3
* Model generated on Jan 31, 2004
* Model format: PSpice
* Darlington macro model
* External node designations
* Node 1 -> Collect
* Node 2 -> Base
* Node 3 -> Emitter
Q1 1 2 4 qmodel
Q2 1 4 3 q1model 11.3767
D1 3 1 dmodel
R1 2 4 10000
R2 4 3 1000
* Default values used in dmodel
*   EG=1.11 TT=0 BV=infinite
.MODEL dmodel d
+IS=1e-12 RS=9.92671 N=0.999184 XTI=2.99919
+CJO=0 VJ=0.75 M=0.33 FC=0.5
.MODEL qmodel npn
+IS=9.95227e-13 BF=123.448 NF=1.11551 VAF=79.7055
+IKF=0.190851 ISE=1.61626e-12 NE=1.58879 BR=0.999157
+NR=0.998586 VAR=92.9909 IKR=0.0999918 ISC=1e-13
+NC=1.99919 RB=9.94154 IRB=0.199184 RBM=9.94149
+RE=0.103128 RC=0.996543 XTB=0.4969 XTI=2.99924 EG=1.11167
+CJE=2.01194e-10 VJE=0.95 MJE=0.23 TF=1e-09
+XTF=1 VTF=10 ITF=0.01 CJC=1.56414e-10
+VJC=0.853057 MJC=0.23 XCJC=0.9 FC=0.5
+TR=1e-07 PTF=0 KF=0 AF=1
.MODEL q1model npn
+IS=9.95227e-13 BF=123.448 NF=1.11551 VAF=79.7055
+IKF=0.190851 ISE=1.61626e-12 NE=1.58879 BR=0.999157
+NR=0.998586 VAR=92.9909 IKR=0.0999918 ISC=1e-13
+NC=1.99919 RB=9.94154 IRB=0.199184 RBM=9.94149
+RE=0.103128 RC=0.996543 XTB=0.4969 XTI=2.99924 EG=1.11167
+CJE=2.01194e-10 VJE=0.95 MJE=0.23 TF=1e-09
+XTF=1 VTF=10 ITF=0.01 CJC=0
+VJC=0.853057 MJC=0.23 XCJC=0.9 FC=0.5
+TR=1e-07 PTF=0 KF=0 AF=1
.ENDS
*******************************************************************
.SUBCKT BDX33C 1 2 3
* Model generated on Dec 24, 2003
* Model format: PSpice
* Darlington macro model
* External node designations
* Node 1 -> Collect
* Node 2 -> Base
* Node 3 -> Emitter
Q1 1 2 4 qmodel
Q2 1 4 3 q1model 11.3524
D1 3 1 dmodel
R1 2 4 10000
R2 4 3 1000
* Default values used in dmodel
*   EG=1.11 TT=0 BV=infinite
.MODEL dmodel d
+IS=1e-12 RS=9.92679 N=0.999268 XTI=2.99927
+CJO=0 VJ=0.75 M=0.33 FC=0.5
.MODEL qmodel npn
+IS=9.96517e-13 BF=123.706 NF=1.08765 VAF=79.7173
+IKF=0.122027 ISE=1.60579e-12 NE=1.58945 BR=0.999264
+NR=0.999167 VAR=92.9992 IKR=0.0999927 ISC=1e-13
+NC=1.99927 RB=9.94157 IRB=0.199268 RBM=9.94157
+RE=0.100179 RC=0.996631 XTB=0.49703 XTI=2.99932 EG=1.11145
+CJE=2.01225e-10 VJE=0.95 MJE=0.23 TF=1e-09
+XTF=1 VTF=10 ITF=0.01 CJC=1.56414e-10
+VJC=0.853047 MJC=0.23 XCJC=0.9 FC=0.5
+TR=1e-07 PTF=0 KF=0 AF=1
.MODEL q1model npn
+IS=9.96517e-13 BF=123.706 NF=1.08765 VAF=79.7173
+IKF=0.122027 ISE=1.60579e-12 NE=1.58945 BR=0.999264
+NR=0.999167 VAR=92.9992 IKR=0.0999927 ISC=1e-13
+NC=1.99927 RB=9.94157 IRB=0.199268 RBM=9.94157
+RE=0.100179 RC=0.996631 XTB=0.49703 XTI=2.99932 EG=1.11145
+CJE=2.01225e-10 VJE=0.95 MJE=0.23 TF=1e-09
+XTF=1 VTF=10 ITF=0.01 CJC=0
+VJC=0.853047 MJC=0.23 XCJC=0.9 FC=0.5
+TR=1e-07 PTF=0 KF=0 AF=1
.ENDS
*******************************************************************
.SUBCKT BDX34B 1 2 3
* Model generated on Jan 31, 2004
* Model format: PSpice
* Darlington macro model
* External node designations
* Node 1 -> Collect
* Node 2 -> Base
* Node 3 -> Emitter
Q1 1 2 4 qmodel
Q2 1 4 3 q1model 11.5248
D1 1 3 dmodel
R1 2 4 10000
R2 4 3 1000
* Default values used in dmodel
*   EG=1.11 TT=0 BV=infinite
.MODEL dmodel d
+IS=1e-12 RS=9.96093 N=0.999455 XTI=2.99945
+CJO=0 VJ=0.75 M=0.33 FC=0.5
.MODEL qmodel pnp
+IS=9.95415e-13 BF=129.468 NF=1.11003 VAF=82.7894
+IKF=0.16855 ISE=1.64286e-12 NE=1.5874 BR=0.999389
+NR=0.998011 VAR=96.4238 IKR=0.0999945 ISC=1e-13
+NC=1.99945 RB=9.97431 IRB=0.199455 RBM=9.97424
+RE=0.103986 RC=0.997005 XTB=0.497049 XTI=2.99952 EG=1.11189
+CJE=1.57148e-10 VJE=2 MJE=2.3e-05 TF=1e-09
+XTF=1 VTF=10 ITF=0.01 CJC=2.46924e-10
+VJC=0.95 MJC=0.244591 XCJC=0.9 FC=0.5
+TR=1e-07 PTF=0 KF=0 AF=1
.MODEL q1model pnp
+IS=9.95415e-13 BF=129.468 NF=1.11003 VAF=82.7894
+IKF=0.16855 ISE=1.64286e-12 NE=1.5874 BR=0.999389
+NR=0.998011 VAR=96.4238 IKR=0.0999945 ISC=1e-13
+NC=1.99945 RB=9.97431 IRB=0.199455 RBM=9.97424
+RE=0.103986 RC=0.997005 XTB=0.497049 XTI=2.99952 EG=1.11189
+CJE=1.57148e-10 VJE=2 MJE=2.3e-05 TF=1e-09
+XTF=1 VTF=10 ITF=0.01 CJC=0
+VJC=0.95 MJC=0.244591 XCJC=0.9 FC=0.5
+TR=1e-07 PTF=0 KF=0 AF=1
.ENDS
*******************************************************************
.SUBCKT BDX34C 1 2 3
* Model generated on Dec 24, 2003
* Model format: PSpice
* Darlington macro model
* External node designations
* Node 1 -> Collect
* Node 2 -> Base
* Node 3 -> Emitter
Q1 1 2 4 qmodel
Q2 1 4 3 q1model 11.5242
D1 1 3 dmodel
R1 2 4 10000
R2 4 3 1000
* Default values used in dmodel
*   EG=1.11 TT=0 BV=infinite
.MODEL dmodel d
+IS=1e-12 RS=9.96109 N=0.999611 XTI=2.99961
+CJO=0 VJ=0.75 M=0.33 FC=0.5
.MODEL qmodel pnp
+IS=9.96197e-13 BF=130.6 NF=1.09163 VAF=82.8066
+IKF=0.124415 ISE=1.63236e-12 NE=1.58838 BR=0.999604
+NR=0.999458 VAR=96.4393 IKR=0.0999961 ISC=1e-13
+NC=1.99961 RB=9.97438 IRB=0.199611 RBM=9.97438
+RE=0.100174 RC=0.996978 XTB=0.497241 XTI=2.99967 EG=1.11187
+CJE=1.57143e-10 VJE=2 MJE=2.3e-05 TF=1e-09
+XTF=1 VTF=10 ITF=0.01 CJC=2.46924e-10
+VJC=0.95 MJC=0.244591 XCJC=0.9 FC=0.5
+TR=1e-07 PTF=0 KF=0 AF=1
.MODEL q1model pnp
+IS=9.96197e-13 BF=130.6 NF=1.09163 VAF=82.8066
+IKF=0.124415 ISE=1.63236e-12 NE=1.58838 BR=0.999604
+NR=0.999458 VAR=96.4393 IKR=0.0999961 ISC=1e-13
+NC=1.99961 RB=9.97438 IRB=0.199611 RBM=9.97438
+RE=0.100174 RC=0.996978 XTB=0.497241 XTI=2.99967 EG=1.11187
+CJE=1.57143e-10 VJE=2 MJE=2.3e-05 TF=1e-09
+XTF=1 VTF=10 ITF=0.01 CJC=0
+VJC=0.95 MJC=0.244591 XCJC=0.9 FC=0.5
+TR=1e-07 PTF=0 KF=0 AF=1
.ENDS
*******************************************************************
*******************************************************************
.SUBCKT BDX53B 1 2 3
* Model generated on Jan 31, 2004
* Model format: PSpice
* Darlington macro model
* External node designations
* Node 1 -> Collect
* Node 2 -> Base
* Node 3 -> Emitter
Q1 1 2 4 qmodel
Q2 1 4 3 q1model 11.9456
D1 3 1 dmodel
R1 2 4 8000
R2 4 3 120
* Default values used in dmodel
*   EG=1.11 TT=0 BV=infinite
.MODEL dmodel d
+IS=1e-12 RS=10 N=1 XTI=3
+CJO=0 VJ=0.75 M=0.33 FC=0.5
.MODEL qmodel npn
+IS=9.87016e-13 BF=153.403 NF=1.2 VAF=78.081
+IKF=0.133947 ISE=1.5267e-12 NE=1.63245 BR=0.999743
+NR=0.994023 VAR=100.425 IKR=0.0999994 ISC=1e-13
+NC=2 RB=10.1734 IRB=0.200041 RBM=10.025
+RE=0.1008 RC=0.997883 XTB=0.496482 XTI=3.00014 EG=1.11532
+CJE=2.58791e-10 VJE=0.95 MJE=0.23 TF=1e-09
+XTF=1 VTF=10 ITF=0.01 CJC=1.54981e-10
+VJC=0.878246 MJC=0.23 XCJC=0.9 FC=0.5
+TR=1e-07 PTF=0 KF=0 AF=1
.MODEL q1model npn
+IS=9.87016e-13 BF=153.403 NF=1.2 VAF=78.081
+IKF=0.133947 ISE=1.5267e-12 NE=1.63245 BR=0.999743
+NR=0.994023 VAR=100.425 IKR=0.0999994 ISC=1e-13
+NC=2 RB=10.1734 IRB=0.200041 RBM=10.025
+RE=0.1008 RC=0.997883 XTB=0.496482 XTI=3.00014 EG=1.11532
+CJE=2.58791e-10 VJE=0.95 MJE=0.23 TF=1e-09
+XTF=1 VTF=10 ITF=0.01 CJC=0
+VJC=0.878246 MJC=0.23 XCJC=0.9 FC=0.5
+TR=1e-07 PTF=0 KF=0 AF=1
.ENDS
*******************************************************************
.SUBCKT BDX53C 1 2 3
* Model generated on Jan 31, 2004
* Model format: PSpice
* Darlington macro model
* External node designations
* Node 1 -> Collect
* Node 2 -> Base
* Node 3 -> Emitter
Q1 1 2 4 qmodel
Q2 1 4 3 q1model 8.40161
D1 3 1 dmodel
R1 2 4 8000
R2 4 3 120
* Default values used in dmodel
*   EG=1.11 TT=0 BV=infinite
.MODEL dmodel d
+IS=1e-12 RS=10 N=1 XTI=3
+CJO=0 VJ=0.75 M=0.33 FC=0.5
.MODEL qmodel npn
+IS=1.20104e-12 BF=160.613 NF=1.2 VAF=78.0305
+IKF=0.154486 ISE=2.74105e-12 NE=1.68339 BR=0.997613
+NR=0.944651 VAR=100.59 IKR=0.0999892 ISC=1e-13
+NC=2 RB=11.2499 IRB=0.211062 RBM=10.1889
+RE=0.223578 RC=1.11789 XTB=0.495729 XTI=2.99866 EG=1.05806
+CJE=2.58424e-10 VJE=0.95 MJE=0.23 TF=1e-09
+XTF=1 VTF=10 ITF=0.01 CJC=1.54982e-10
+VJC=0.878229 MJC=0.23 XCJC=0.9 FC=0.5
+TR=1e-07 PTF=0 KF=0 AF=1
.MODEL q1model npn
+IS=1.20104e-12 BF=160.613 NF=1.2 VAF=78.0305
+IKF=0.154486 ISE=2.74105e-12 NE=1.68339 BR=0.997613
+NR=0.944651 VAR=100.59 IKR=0.0999892 ISC=1e-13
+NC=2 RB=11.2499 IRB=0.211062 RBM=10.1889
+RE=0.223578 RC=1.11789 XTB=0.495729 XTI=2.99866 EG=1.05806
+CJE=2.58424e-10 VJE=0.95 MJE=0.23 TF=1e-09
+XTF=1 VTF=10 ITF=0.01 CJC=0
+VJC=0.878229 MJC=0.23 XCJC=0.9 FC=0.5
+TR=1e-07 PTF=0 KF=0 AF=1
.ENDS
*******************************************************************
.SUBCKT BDX54B 1 2 3
* Model generated on Jan 31, 2004
* Model format: PSpice
* Darlington macro model
* External node designations
* Node 1 -> Collect
* Node 2 -> Base
* Node 3 -> Emitter
Q1 1 2 4 qmodel
Q2 1 4 3 q1model 8.33943
D1 1 3 dmodel
R1 2 4 8000
R2 4 3 120
* Default values used in dmodel
*   EG=1.11 TT=0 BV=infinite
.MODEL dmodel d
+IS=1e-12 RS=10 N=1 XTI=3
+CJO=0 VJ=0.75 M=0.33 FC=0.5
.MODEL qmodel pnp
+IS=1.4554e-12 BF=188.357 NF=1.2 VAF=105.353
+IKF=0.124891 ISE=3.85559e-13 NE=1.51221 BR=0.996693
+NR=0.914215 VAR=101.606 IKR=0.0999754 ISC=1e-13
+NC=2 RB=13.4247 IRB=0.231 RBM=10.9398
+RE=0.107708 RC=1.10559 XTB=0.488759 XTI=2.99693 EG=1.05
+CJE=2.6466e-10 VJE=0.95 MJE=0.23 TF=1e-09
+XTF=1 VTF=10 ITF=0.01 CJC=2.49703e-10
+VJC=0.81223 MJC=0.23 XCJC=0.9 FC=0.5
+TR=1e-07 PTF=0 KF=0 AF=1
.MODEL q1model pnp
+IS=1.4554e-12 BF=188.357 NF=1.2 VAF=105.353
+IKF=0.124891 ISE=3.85559e-13 NE=1.51221 BR=0.996693
+NR=0.914215 VAR=101.606 IKR=0.0999754 ISC=1e-13
+NC=2 RB=13.4247 IRB=0.231 RBM=10.9398
+RE=0.107708 RC=1.10559 XTB=0.488759 XTI=2.99693 EG=1.05
+CJE=2.6466e-10 VJE=0.95 MJE=0.23 TF=1e-09
+XTF=1 VTF=10 ITF=0.01 CJC=0
+VJC=0.81223 MJC=0.23 XCJC=0.9 FC=0.5
+TR=1e-07 PTF=0 KF=0 AF=1
.ENDS
*******************************************************************
.SUBCKT BDX54C 1 2 3
* Model generated on Jan 31, 2004
* Model format: PSpice
* Darlington macro model
* External node designations
* Node 1 -> Collect
* Node 2 -> Base
* Node 3 -> Emitter
Q1 1 2 4 qmodel
Q2 1 4 3 q1model 8.33905
D1 1 3 dmodel
R1 2 4 8000
R2 4 3 120
* Default values used in dmodel
*   EG=1.11 TT=0 BV=infinite
.MODEL dmodel d
+IS=1e-12 RS=10 N=1 XTI=3
+CJO=0 VJ=0.75 M=0.33 FC=0.5
.MODEL qmodel pnp
+IS=1.56186e-12 BF=188.227 NF=1.1739 VAF=105.358
+IKF=0.113314 ISE=3.87694e-13 NE=1.50183 BR=0.996711
+NR=0.914768 VAR=101.604 IKR=0.0999754 ISC=1e-13
+NC=2 RB=13.4402 IRB=0.231192 RBM=10.9425
+RE=0.113908 RC=1.10586 XTB=0.488781 XTI=2.99692 EG=1.05
+CJE=2.60341e-10 VJE=0.95 MJE=0.23 TF=1e-09
+XTF=1 VTF=10 ITF=0.01 CJC=2.47462e-10
+VJC=0.95 MJC=0.23 XCJC=0.9 FC=0.5
+TR=1e-07 PTF=0 KF=0 AF=1
.MODEL q1model pnp
+IS=1.56186e-12 BF=188.227 NF=1.1739 VAF=105.358
+IKF=0.113314 ISE=3.87694e-13 NE=1.50183 BR=0.996711
+NR=0.914768 VAR=101.604 IKR=0.0999754 ISC=1e-13
+NC=2 RB=13.4402 IRB=0.231192 RBM=10.9425
+RE=0.113908 RC=1.10586 XTB=0.488781 XTI=2.99692 EG=1.05
+CJE=2.60341e-10 VJE=0.95 MJE=0.23 TF=1e-09
+XTF=1 VTF=10 ITF=0.01 CJC=0
+VJC=0.95 MJC=0.23 XCJC=0.9 FC=0.5
+TR=1e-07 PTF=0 KF=0 AF=1
.ENDS
*******************************************************************
*******************************************************************
.SUBCKT TIP122 1 2 3
* Model generated on Dec 19, 2003
* Model format: PSpice
* Darlington macro model
* External node designations
* Node 1 -> Collect
* Node 2 -> Base
* Node 3 -> Emitter
Q1 1 2 4 qmodel
Q2 1 4 3 q1model 2.7545
D1 3 1 dmodel
R1 2 4 10000
R2 4 3 1000
* Default values used in dmodel
*   EG=1.11 TT=0 BV=infinite
.MODEL dmodel d
+IS=1e-12 RS=10 N=1 XTI=3
+CJO=0 VJ=0.75 M=0.33 FC=0.5
.MODEL qmodel npn
+IS=1.15528e-13 BF=387.828 NF=0.937439 VAF=30
+IKF=0.270029 ISE=5.36359e-11 NE=1.54544 BR=0.1
+NR=1.5 VAR=134.979 IKR=0.109764 ISC=1.00329e-13
+NC=1.97549 RB=4.9473 IRB=0.200762 RBM=4.9473
+RE=0.0964614 RC=0.482307 XTB=0.580269 XTI=2.92642 EG=1.05
+CJE=2.08206e-10 VJE=0.945586 MJE=0.23 TF=1e-09
+XTF=1 VTF=10 ITF=0.01 CJC=1.67927e-10
+VJC=0.754327 MJC=0.289398 XCJC=0.9 FC=0.5
+TR=1e-07 PTF=0 KF=0 AF=1
.MODEL q1model npn
+IS=1.15528e-13 BF=387.828 NF=0.937439 VAF=30
+IKF=0.270029 ISE=5.36359e-11 NE=1.54544 BR=0.1
+NR=1.5 VAR=134.979 IKR=0.109764 ISC=1.00329e-13
+NC=1.97549 RB=4.9473 IRB=0.200762 RBM=4.9473
+RE=0.0964614 RC=0.482307 XTB=0.580269 XTI=2.92642 EG=1.05
+CJE=2.08206e-10 VJE=0.945586 MJE=0.23 TF=1e-09
+XTF=1 VTF=10 ITF=0.01 CJC=0
+VJC=0.754327 MJC=0.289398 XCJC=0.9 FC=0.5
+TR=1e-07 PTF=0 KF=0 AF=1
.ENDS
*******************************************************************
.SUBCKT TIP127 1 2 3
* Model generated on Dec 26, 2003
* Model format: PSpice
* Darlington macro model
* External node designations
* Node 1 -> Collect
* Node 2 -> Base
* Node 3 -> Emitter
Q1 1 2 4 qmodel
Q2 1 4 3 q1model 2.84905
D1 1 3 dmodel
R1 2 4 10000
R2 4 3 1000
* Default values used in dmodel
*   EG=1.11 TT=0 BV=infinite
.MODEL dmodel d
+IS=1e-12 RS=10 N=1 XTI=3
+CJO=0 VJ=0.75 M=0.33 FC=0.5
.MODEL qmodel pnp
+IS=2.2383e-14 BF=390.271 NF=0.874443 VAF=38.5083
+IKF=0.202108 ISE=1.49947e-10 NE=1.64874 BR=0.1
+NR=1.32278 VAR=134.629 IKR=0.177707 ISC=1.03339e-13
+NC=1.97553 RB=4.89811 IRB=0.200734 RBM=4.89811
+RE=0.089979 RC=0.449895 XTB=0.584937 XTI=2.92881 EG=1.05
+CJE=2.09764e-10 VJE=0.95 MJE=0.23 TF=1e-09
+XTF=1 VTF=10 ITF=0.01 CJC=1.53285e-10
+VJC=0.95 MJC=0.23 XCJC=0.9 FC=0.5
+TR=1e-07 PTF=0 KF=0 AF=1
.MODEL q1model pnp
+IS=2.2383e-14 BF=390.271 NF=0.874443 VAF=38.5083
+IKF=0.202108 ISE=1.49947e-10 NE=1.64874 BR=0.1
+NR=1.32278 VAR=134.629 IKR=0.177707 ISC=1.03339e-13
+NC=1.97553 RB=4.89811 IRB=0.200734 RBM=4.89811
+RE=0.089979 RC=0.449895 XTB=0.584937 XTI=2.92881 EG=1.05
+CJE=2.09764e-10 VJE=0.95 MJE=0.23 TF=1e-09
+XTF=1 VTF=10 ITF=0.01 CJC=0
+VJC=0.95 MJC=0.23 XCJC=0.9 FC=0.5
+TR=1e-07 PTF=0 KF=0 AF=1
.ENDS
*******************************************************************
*TIP141 MCE Nodes: C B E 7/6/95
*MCE  80V  10A
.SUBCKT XTIP141   1 2 3
Q1 1 2 4 QPWR .1
Q2 1 4 3 QPWR
R1 2 4  8K
R2 4 3  40
D1 3 1  DSUB
.MODEL QPWR NPN(IS=12P NF=1 BF=99.9 VAF=161 IKF=8 ISE=981P NE=2
+ BR=4 NR=1 VAR=20 IKR=12 RE=40M RB=.16 RC=16M XTB=1.5
+ CJE=1.34N VJE=.74 MJE=.45 CJC=193P VJC=1.1 MJC=.24 TF=98.5N TR=4.25U)
.MODEL DSUB D(IS=12P N=1 RS=40M BV=80 IBV=.001 CJO=193P TT=4.25U)
.ENDS XTIP141
********************************************************************
.SUBCKT BD681 1 2 3
* Model generated on Feb 28, 2004
* Model format: PSpice
* Darlington macro model
* External node designations
* Node 1 -> Collect
* Node 2 -> Base
* Node 3 -> Emitter
Q1 1 2 4 qmodel
Q2 1 4 3 q1model 5.21716
D1 3 1 dmodel
R1 2 4 8000
R2 4 3 120
* Default values used in dmodel
*   EG=1.11 TT=0 BV=infinite
.MODEL dmodel d
+IS=1e-12 RS=9.53186 N=0.964987 XTI=2.96499
+CJO=0 VJ=0.75 M=0.33 FC=0.5
.MODEL qmodel npn
+IS=6.82736e-17 BF=43.4441 NF=0.85 VAF=30
+IKF=1.14362 ISE=9.48937e-15 NE=2.04295 BR=0.665831
+NR=1.5 VAR=64.8234 IKR=0.0980345 ISC=9.48937e-15
+NC=1 RB=20.4512 IRB=0.277791 RBM=16.9143
+RE=0.574152 RC=6.88011 XTB=0.401039 XTI=2.96301 EG=1.05
+CJE=1e-11 VJE=0.75 MJE=0.33 TF=1e-09
+XTF=1 VTF=10 ITF=0.01 CJC=1e-11
+VJC=0.75 MJC=0.33 XCJC=0.9 FC=0.5
+TR=1e-07 PTF=0 KF=0 AF=1
.MODEL q1model npn
+IS=6.82736e-17 BF=43.4441 NF=0.85 VAF=30
+IKF=1.14362 ISE=9.48937e-15 NE=2.04295 BR=0.665831
+NR=1.5 VAR=64.8234 IKR=0.0980345 ISC=9.48937e-15
+NC=1 RB=20.4512 IRB=0.277791 RBM=16.9143
+RE=0.574152 RC=6.88011 XTB=0.401039 XTI=2.96301 EG=1.05
+CJE=1e-11 VJE=0.75 MJE=0.33 TF=1e-09
+XTF=1 VTF=10 ITF=0.01 CJC=0
+VJC=0.75 MJC=0.33 XCJC=0.9 FC=0.5
+TR=1e-07 PTF=0 KF=0 AF=1
.ENDS
********************************************************************
.SUBCKT BD682 1 2 3
* Model generated on Feb 28, 2004
* Model format: PSpice
* Darlington macro model
* External node designations
* Node 1 -> Collect
* Node 2 -> Base
* Node 3 -> Emitter
Q1 1 2 4 qmodel
Q2 1 4 3 q1model 2.46191
D1 1 3 dmodel
R1 2 4 8000
R2 4 3 120
* Default values used in dmodel
*   EG=1.11 TT=0 BV=infinite
.MODEL dmodel d
+IS=1e-12 RS=10 N=1 XTI=3
+CJO=0 VJ=0.75 M=0.33 FC=0.5
.MODEL qmodel pnp
+IS=2.23835e-12 BF=149.682 NF=1.2 VAF=59.0895
+IKF=0.118079 ISE=9.09119e-14 NE=1.42175 BR=0.587475
+NR=0.75 VAR=100.388 IKR=0.0934405 ISC=9.09118e-14
+NC=2 RB=15.5445 IRB=0.450416 RBM=12.8364
+RE=0.0939759 RC=2.76027 XTB=0.497353 XTI=2.9942 EG=1.05
+CJE=1e-11 VJE=0.75 MJE=0.33 TF=1e-09
+XTF=1 VTF=10 ITF=0.01 CJC=1e-11
+VJC=0.75 MJC=0.33 XCJC=0.9 FC=0.5
+TR=1e-07 PTF=0 KF=0 AF=1
.MODEL q1model pnp
+IS=2.23835e-12 BF=149.682 NF=1.2 VAF=59.0895
+IKF=0.118079 ISE=9.09119e-14 NE=1.42175 BR=0.587475
+NR=0.75 VAR=100.388 IKR=0.0934405 ISC=9.09118e-14
+NC=2 RB=15.5445 IRB=0.450416 RBM=12.8364
+RE=0.0939759 RC=2.76027 XTB=0.497353 XTI=2.9942 EG=1.05
+CJE=1e-11 VJE=0.75 MJE=0.33 TF=1e-09
+XTF=1 VTF=10 ITF=0.01 CJC=0
+VJC=0.75 MJC=0.33 XCJC=0.9 FC=0.5
+TR=1e-07 PTF=0 KF=0 AF=1
.ENDS




