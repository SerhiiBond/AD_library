*SI3442DV  MCE  5-27-97
*20V 4A 0.065ohm Power MOSFET pkg:TSOP-6 1,3,4
.SUBCKT SI3442DV 10 20 40 40
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  29.9M
RS  40  3  2.62M
RG  20  2  37.5
CGS  2  3  420P
EGD 12  0  2  1  1
VFB 14  0  0
FFB  2  1  VFB  1
CGD 13 14  317P
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD  3 10  DSUB
LS  30 40  7.5N
.MODEL DMOS NMOS (LEVEL=3 VMAX=41.7K THETA=80M ETA=2M VTO=0.6 KP=79.4)
.MODEL DCGD D (CJO=317P VJ=0.6 M=0.68)
.MODEL DSUB D (IS=16.6N N=1.5 RS=0 BV=20 CJO=352P VJ=0.8 M=0.42 TT=40N)
.MODEL DLIM D (IS=100U)
.ENDS 