*DZ23C12 MCE 4/9/98
*Ref: Diodes Incorporated, 1994
*12V 350mW Si Dual Zener pkg:TO236AA 1,3,2
.SUBCKT DZ23C12 1 2 3
*      TERMINALS A K A
XA 1 2 DDZ23C12
XB 3 2 DDZ23C12
.ENDS DZ23C12


.SUBCKT DDZ23C12  1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  11.46
.MODEL DF D (IS=1.76N RS=0.12 N=1.7 CJO=42.7P VJ=1 M=0.33 TT=50.1N)
.MODEL DR D (IS=16.5U RS=7.5 N=3.4)
.ENDS DDZ23C12