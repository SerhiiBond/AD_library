*SI4480DY  MCE  5-27-97
*80V 6A 0.028ohm Power MOSFET pkg:SMD8A 8,4,1
.SUBCKT SI4480DY 10 20 40 40
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  12.3M
RS  40  3  1.7M
RG  20  2  25
CGS  2  3  1.81N
EGD 12  0  2  1  1
VFB 14  0  0
FFB  2  1  VFB  1
CGD 13 14  1.3N
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD  3 10  DSUB
LS  30 40  7.5N
.MODEL DMOS NMOS (LEVEL=3 VMAX=167K THETA=80M ETA=2M VTO=2 KP=131)
.MODEL DCGD D (CJO=1.3N VJ=0.6 M=0.68)
.MODEL DSUB D (IS=24.9N N=1.5 RS=41.7M BV=80 CJO=927P VJ=0.8 M=0.42 TT=50N)
.MODEL DLIM D (IS=100U)
.ENDS 