*                D G S
.SUBCKT ZVP4424A 3 4 5
M1 3 2 5 5 P4424AM
RG 4 2 140
RL 3 5 4E9
D1 3 5 P4424AD
.MODEL P4424AM PMOS VTO=-1.5 RS=1.245 RD=6.2 IS=1E-15 KP=0.52
+CGSO=98.8E-12 CGDO=3.2E-12 CBD=65.3E-12 PB=1
.MODEL P4424AD D IS=9.36E-13 RS=.196 N=1.045
.ENDS ZVP4424A
