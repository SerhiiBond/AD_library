*SI4925DY  MCE  5-28-97
* jjt 4/4/2002: changed VTO to -1V to match  S-51642�Rev. C, 17-Mar-97 datasheet
*30V 6A 0.031ohm Dual Power MOSFET pkg:SMD8A (A:8,2,1)(B:6,4,3)
.SUBCKT SI4925DY 10 20 40 40
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  13.7M
RS  40  3  1.78M
RG  20  2  24.6
CGS  2  3  1.79N
EGD 12  0  1  2  1
VFB 14  0  0
FFB  1  2  VFB  1
CGD 13 14  2.07N
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD 10  3  DSUB
LS  30 40  7.5N
.MODEL DMOS PMOS (LEVEL=3 VMAX=62.5K THETA=80M ETA=2M VTO=-1 KP=81.4)
.MODEL DCGD D (CJO=2.07N VJ=0.6 M=0.68)
.MODEL DSUB D (IS=25.3N N=1.5 RS=65.6M BV=30 CJO=2.26N VJ=0.8 M=0.42 TT=50N)
.MODEL DLIM D (IS=100U)
.ENDS 