*SI6332DQ  MCE  5-28-97
* jjt 4/4/2002: changed sign of VTO to match S-49520-Rev. C,18-Dec-96 datasheet
*30V 4A 0.037ohm Triple Power MOSFET pkg:SMD28 (A:1,4,26)(B:6,9,21)(C:11,14,16)
.SUBCKT SI6332DQ 10 20 40 40
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  16.6M
RS  40  3  1.93M
RG  20  2  33.3
CGS  2  3  1.16N
EGD 12  0  1  2  1
VFB 14  0  0
FFB  1  2  VFB  1
CGD 13 14  1.55N
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD 10  3  DSUB
LS  30 40  7.5N
.MODEL DMOS PMOS (LEVEL=3 VMAX=62.5K THETA=80M ETA=2M VTO=-1 KP=34.9)
.MODEL DCGD D (CJO=1.55N VJ=0.6 M=0.68)
.MODEL DSUB D (IS=18.7N N=1.5 RS=11.1M BV=30 CJO=904P VJ=0.8 M=0.42 TT=50N)
.MODEL DLIM D (IS=100U)
.ENDS 