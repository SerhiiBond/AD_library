*SI6933DQ  MCE  5-28-97
*30V 4A 0.059ohm Dual Power MOSFET pkg:SMD8B (A:1,4,3)(B:8,5,6)
.SUBCKT SI6933DQ 10 20 40 40
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  27M
RS  40  3  2.48M
RG  20  2  42.9
CGS  2  3  1.07N
EGD 12  0  1  2  1
VFB 14  0  0
FFB  1  2  VFB  1
CGD 13 14  1.03N
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD 10  3  DSUB
LS  30 40  7.5N
.MODEL DMOS PMOS (LEVEL=3 VMAX=62.5K THETA=80M ETA=2M VTO=-1 KP=28.7)
.MODEL DCGD D (CJO=1.03N VJ=0.6 M=0.68)
.MODEL DSUB D (IS=14.5N N=1.5 RS=5.71M BV=30 CJO=471P VJ=0.8 M=0.42 TT=30N)
.MODEL DLIM D (IS=100U)
.ENDS 