*FDV302P at Temp. Electrical Model 
*-------------------------------------
.SUBCKT FDV302P 20 10 30
*20=DRAIN 10=GATE 30=SOURCE 50=VTEMP
Rg 10 11x 1
Rdu 12x 1 1u
M1 2 1 4x 4x DMOS L=1u W=1u
.MODEL DMOS PMOS(VTO=-0.83 KP=1.53E-1
+THETA=0.25 VMAX=2E5 LEVEL=3)
Cgs 1 5x 32p
Rd 20 4 1.4
Dds 4 5x DDS
.MODEL DDS D(M=2.91E-1 VJ=4.64E-1 CJO=14.1p)
Dbody 20 5x DBODY
.MODEL DBODY D(IS=7.94E-8 N=2.460181 RS=.021333 TT=52.03n)
Ra 4 2 1.4 
Rs 5x 5 0.5m
Ls 5 30 0.5n
M2 1 8 6 6 INTER
E2 8 6 4 1 2
.MODEL INTER PMOS(VTO=0 KP=10 LEVEL=1)
Cgdmax 7 4 35.6p
Rcgd 7 4 10meg
Dgd 4 6 DGD
Rdgd 4 6 10meg
.MODEL DGD D(M=5.5E-1 VJ=2.6E-3 CJO=35.6p)
M3 7 9 1 1 INTER
E3 9 1 4 1 -2
*ZX SECTION
EOUT 4x 6x poly(2) (1x,0) (3x,0) 0 0 0 0 1
FCOPY 0 3x VSENSE 1
RIN 1x 0 1G
VSENSE 6x 5x 0
RREF 3x 0 10m
*TEMP SECTION
*ED 101 0 VALUE {V(50,100)}
VAMB 100 0 25
EKP 1x 0 101 0 2.9
*VTO TEMP SECTION
EVTO 102 0 101 0 .0016
EVT 11x 12x 102 0 1
*DIODE THEMO BREAKDOWN SECTION
EBL VB1 VB2 101 0 .08
VBLK VB2 0 25
D DB1 20 DBLK
.MODEL DBLK D(IS=1E-14 CJO=.1p RS=.1)
EDB 0 DB1 VB1 0 1
.ENDS FDV302P
*FDV302P (Rev.B) 10/23/01 **ST

