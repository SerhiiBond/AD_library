*DL4755A MCE 4/8/98
*Ref: Diodes Incorporated, 1994
*43V 1W Si Zener pkg:DL-41 1,2
.SUBCKT DL4755A  1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  42.32
.MODEL DF D (IS=5.02N RS=42M N=1.7 CJO=37.1P VJ=1 M=0.33 TT=50.1N)
.MODEL DR D (IS=1.1M RS=21 N=11)
.ENDS