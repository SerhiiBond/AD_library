*Si4412DY Siliconix 2-Oct-96
*N-Channel DMOS Subcircuit Model
.SUBCKT Si4412DY 4 1 2 2
M1 3 1 2 2 NMOS W=1755000U L=0.5U
R1 4 3 RTEMP 135E-4
CGS 1 2 550PF
CGD 1 6 550PF
DMIN 6 4 DMIN
DMAX 6 1 DMAX
DBODY 2 4 DBODY
.MODEL NMOS NMOS(LEVEL=3 TOX=5.00E-8 RS=45.5E-4 RD=0 LD=0
+ NSUB=1.85E+17 UO=400 VMAX=0 ETA=3.0E-4 XJ=5E-7
+ KAPPA=0.25 CGBO=0 TPG=1 DELTA=0.1 CGSO=0 CGDO=0
+ IS=0 KP=1.5E-5 NFS=.1E+12)
.MODEL DMIN D(CJO=530E-12 VJ=0.15 M=0.5 FC=0.5 IS=1E-20)
.MODEL DMAX D(CJO=650E-12 VJ=0.6 M=0.45 FC=0.5 IS=1E-22)
.MODEL DBODY D(CJO=950E-12 VJ=0.8 M=0.36 FC=0.5 N=1 IS=1E-15
+ TT=1.4E-8 BV=40)
.MODEL RTEMP R(TC1=4E-3 TC2=12E-6)
.ENDS 