*BZT52C8V2 MCE 4/8/98
*Ref: Diodes Incorporated, 1994
*8.2V 410mW Si Zener pkg:60A2 1,2
.SUBCKT BZT52C8V2 1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  7.678
.MODEL DF D (IS=2.06N RS=0.102 N=1.7 CJO=38.1P VJ=0.75 M=0.33 TT=50.1N)
.MODEL DR D (IS=365N RS=4.5 N=2)
.ENDS