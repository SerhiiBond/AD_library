*IRFK3D450 MCE  12/12/97
*Ref: International Rectifier Product Digest '94
*500V 33A .0364ohm Power MOSFET pkg:TO-126 2,3,1
*SYM=POWMOSN
*pn,29/06/2000,merged both parts into 1 subckt

.SUBCKT IRFK3D450 D1 G1 S1D2 G2 S2
X1 D1 G1 S1D2 MIRFK3D450
X2 S1D2 G2 S2 MIRFK3D450
.ENDS

.SUBCKT MIRFK3D450 10 20 40
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  16.3M
RS  40  3  1.91M
RG  20  2  4.55
CGS  2  3  951P
EGD 12  0  2  1  1
VFB 14  0  0
FFB  2  1  VFB  1
CGD 13 14  1.21N
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD  3 10  DSUB
LS  30 40  7.5N
.MODEL DMOS NMOS (LEVEL=3 VMAX=1.04MEG THETA=58.1M ETA=2M VTO=3.1 KP=9.11)
.MODEL DCGD D (CJO=1.21N VJ=0.6 M=0.68)
.MODEL DSUB D (IS=137N N=1.5 RS=18.2M BV=500 IBV=3M CJO=1.84N VJ=0.8 M=0.42 TT=403N)
.MODEL DLIM D (IS=100U)
.ENDS 


