*SiSi3454DV Siliconix 13-Dec-96
*N-Channel DMOS Subcircuit Model
.SUBCKT Si3454DV 4 1 2 2
M1 3 1 2 2 NMOS W=578370U L=0.5U
R1 4 3 RTEMP 36.54M
CGS 1 2 60PF
CGD 1 6 160PF
DMIN 6 4 DMIN
DMAX 6 1 DMAX
DBODY 2 4 DBODY
.MODEL NMOS NMOS(LEVEL=3 TOX=5.00E-8 RS=0.001 RD=0 LD=0
+ NSUB=2.82E+17 VTO=2.963 UO=800 VMAX=0 ETA=3E-4 XJ=0.5E-6
+ KAPPA=0 CGBO=0 TPG=1 DELTA=0.1 CGSO=0 CGDO=0
+ IS=0 KP=9.3913U)
.MODEL DMIN D(CJO=270E-12 VJ=0.09 M=0.54 FC=0.5 IS=1E-21)
.MODEL DMAX D(CJO=270E-12 VJ=0.09 M=0.54 FC=0.5 IS=1E-21)
.MODEL DBODY D(CJO=435E-12 VJ=0.21 M=0.29 FC=0.5 N=1 IS=1E-21
+ TT=1.4E-8 BV=40)
.MODEL RTEMP R(TC1=0.3E-2 TC2=5.0E-6)
.ENDS 