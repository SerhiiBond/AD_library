*SI9424DY  MCE  5-28-97
* jjt 4/4/2002: changed VTO to -0.6V to match S-56950�Rev. E, 11-Jan-99 datasheet
*12V 8A 0.022ohm Power MOSFET pkg:SMD8A 8,4,1
.SUBCKT SI9424DY 10 20 40 40
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  9.45M
RS  40  3  1.55M
RG  20  2  19.5
CGS  2  3  2.6N
EGD 12  0  1  2  1
VFB 14  0  0
FFB  1  2  VFB  1
CGD 13 14  3.57N
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD 10  3  DSUB
LS  30 40  7.5N
.MODEL DMOS PMOS (LEVEL=3 VMAX=25K THETA=80M ETA=2M VTO=-0.6 KP=291)
.MODEL DCGD D (CJO=3.57N VJ=0.6 M=0.68)
.MODEL DSUB D (IS=441N N=1.5 RS=9.35M BV=12 CJO=2.46N VJ=0.8 M=0.42 TT=70N)
.MODEL DLIM D (IS=100U)
.ENDS 