*DZ23C5V1 MCE 4/9/98
*Ref: Diodes Incorporated, 1994
*5.1V 350mW Si Dual Zener pkg:TO236AA 1,3,2
.SUBCKT DZ23C5V1 1 2 3
*      TERMINALS A K A
XA 1 2 DDZ23C5V1
XB 3 2 DDZ23C5V1
.ENDS DZ23C5V1


.SUBCKT DDZ23C5V1 1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  4.492
.MODEL DF D (IS=1.76N RS=0.12 N=1.7 CJO=66.2P VJ=0.75 M=0.33 TT=50.1N)
.MODEL DR D (IS=462U RS=18 N=8.1)
.ENDS DDZ23C5V1