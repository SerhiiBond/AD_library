*BZT52C4V7 MCE 4/8/98
*Ref: Diodes Incorporated, 1994
*4.7V 410mW Si Zener pkg:60A2 1,2
.SUBCKT BZT52C4V7 1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  4.037
.MODEL DF D (IS=2.06N RS=0.102 N=1.7 CJO=87.7P VJ=0.75 M=0.33 TT=50.1N)
.MODEL DR D (IS=838U RS=24 N=11)
.ENDS