*DZ23C3V6 MCE 4/9/98
*Ref: Diodes Incorporated, 1994
*3.6V 350mW Si Dual Zener pkg:TO236AA 1,3,2
.SUBCKT DZ23C3V6 1 2 3
*      TERMINALS A K A
XA 1 2 DDZ23C3V6
XB 3 2 DDZ23C3V6
.ENDS DZ23C3V6


.SUBCKT DDZ23C3V6 1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  2.891
.MODEL DF D (IS=1.76N RS=0.12 N=1.7 CJO=112P VJ=0.75 M=0.33 TT=50.1N)
.MODEL DR D (IS=1.11M RS=28.5 N=13)
.ENDS DDZ23C3V6