*Si9947DY Siliconix 13-Dec-96
*P-Channel DMOS Subcircuit Model
.SUBCKT Si9947DY 4 1 2 2
M1 3 1 2 2 PMOS W=201968U L=0.5U
R1 4 3 RTEMP 25M
CGS 1 2 360PF
CGD 1 6 455PF
DMIN 4 6 DMIN
DMAX 1 6 DMAX
DBODY 4 2 DBODY
.MODEL PMOS PMOS(LEVEL=3 TOX=50N RS=10M RD=0 LD=0
+ NSUB=2.86E+16 VTO=-3.05 UO=250 VMAX=0 ETA=300U XJ=500N THETA=0
+ KAPPA=10M CGBO=0 TPG=-1 DELTA=0 CGSO=0 CGDO=0 IS=0 KP=11.5U)
.MODEL DMIN D(CJO=840P VJ=0.4 M=0.75 FC=0.56 IS=1E-20)
.MODEL DMAX D(CJO=900P VJ=0.5 M=0.5 FC=0.5 IS=1E-22)
.MODEL DBODY D(CJO=1040P VJ=0.09 M=0.25 FC=0.5 N=1 IS=1E-18
+ TT=100N BV=40)
.MODEL RTEMP R(TC1=1.5M TC2=5U)
.ENDS Si9947DY