*SI9803DY  MCE  5-28-97
*20V 6A 0.038ohm Reduced Power MOSFET pkg:SMD8A 8,4,1
.SUBCKT SI9803DY 10 20 40 40
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  17.1M
RS  40  3  1.95M
RG  20  2  25.4
CGS  2  3  1.24N
EGD 12  0  1  2  1
VFB 14  0  0
FFB  1  2  VFB  1
CGD 13 14  5.39N
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD 10  3  DSUB
LS  30 40  7.5N
.MODEL DMOS PMOS (LEVEL=3 VMAX=41.7K THETA=80M ETA=2M VTO=-0.6 KP=137)
.MODEL DCGD D (CJO=5.39N VJ=0.6 M=0.68)
.MODEL DSUB D (IS=24.5N N=1.5 RS=0 BV=20 CJO=1.41N VJ=0.8 M=0.42 TT=80N)
.MODEL DLIM D (IS=100U)
.ENDS 