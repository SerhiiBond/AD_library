*DZ23C16 MCE 4/9/98
*Ref: Diodes Incorporated, 1994
*16V 350mW Si Dual Zener pkg:TO236AA 1,3,2
.SUBCKT DZ23C16 1 2 3
*      TERMINALS A K A
XA 1 2 DDZ23C16
XB 3 2 DDZ23C16
.ENDS DZ23C16


.SUBCKT DDZ23C16  1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  15.44
.MODEL DF D (IS=1.76N RS=0.12 N=1.7 CJO=35.8P VJ=1 M=0.33 TT=50.1N)
.MODEL DR D (IS=141U RS=12 N=5.4)
.ENDS DDZ23C16