*BZT52C5V1 MCE 4/8/98
*Ref: Diodes Incorporated, 1994
*5.1V 410mW Si Zener pkg:60A2 1,2
.SUBCKT BZT52C5V1 1 2
*    TERMINALS:  A K
D1 1 2  DF
DZ 3 1  DR
VZ 2 3  4.492
.MODEL DF D (IS=2.06N RS=0.102 N=1.7 CJO=77.6P VJ=0.75 M=0.33 TT=50.1N)
.MODEL DR D (IS=462U RS=18 N=8.1)
.ENDS